`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// This document contains information prorietary to the CSULB student that created
// the file -  any reuse without adequate approval and documentation is prohibited
//
// File Name: Receive.v
// Project: 3
// Created by <Hung Le> on <April 16, 2019>
// Copright @ 2019 <Hung Le>. All rights reserved
//
// Purpose: This module implements functionality of the receive engine. Control
//	block generates BTU and DONE signals to initiate data collection. They are 
//	generated by control signals from state machine (START,DOIT). Data flow block
//	shifts in data and right justifies it. Then the data is analyzed to ensure the 
// correct parity, correct number of bits, and correct stop bit. Output data of 
// receive is 8-bits. Rxrdy will be set when the engine is ready to sample the 
// next data string. 
//
// In submitting this file for class work at CSULB
// I am confirming that this is my work and the work of no one else. 
// 
// In submitting this code I acknowledge that plagiarism in student project
// work is subject to dismissal from the class. 
//////////////////////////////////////////////////////////////////////////////////
module Receive(clk, rst, k, k_half, eight, pen, ohel, read, RX, rxrdy,
					OVF, FERR, PERR, rx_data);
	input clk, rst, RX, eight, pen, ohel;
	input [7:0] read; 
	input [18:0] k, k_half;
	
	output wire OVF, FERR, PERR, rxrdy;
	output wire [7:0] rx_data;
	assign rx_data = (eight)?	remap_out[7:0] : {1'b0,remap_out[6:0]};
	///////////////////////////////////////////////////////////////////
	//////////////////////RECEIVE ENGINE CONTROL///////////////////////
	///////////////////////////////////////////////////////////////////
	wire SH, DONE, BTU;
	wire [18:0] btu_comp;
	reg  [3:0] 	done_comp, D1, Q1; 
	reg  START, DOIT, nSTART, nDOIT;
	reg  [1:0] NS, PS;
	reg  [18:0] D, Q;
	
	/*****************************************************************/
	//State machine
	/*****************************************************************/
	always @ (posedge clk, posedge rst)
		if(rst)
			{PS,START,DOIT} <= 4'b0;
			
		else
			{PS,START,DOIT} <= {NS,nSTART,nDOIT};
			
	always @ (*) 
		casez({PS, RX, DONE, BTU})
			//state 1 - output: start = 0, doit = 0
			5'b00_1_?_?: {NS,nSTART,nDOIT} = 4'b00_0_0;			
			5'b00_0_?_?: {NS,nSTART,nDOIT} = 4'b01_0_0;
			
			//state 2 - output: start = 1, doit = 1
			5'b01_1_?_?: {NS,nSTART,nDOIT} = 4'b00_1_1;
			5'b01_0_?_0: {NS,nSTART,nDOIT} = 4'b01_1_1;
			5'b01_0_?_1: {NS,nSTART,nDOIT} = 4'b10_1_1;
			
			//state 3 - output: start = 0, doit = 1
			5'b10_?_0_?: {NS,nSTART,nDOIT} = 4'b10_0_1;
			5'b10_?_1_?: {NS,nSTART,nDOIT} = 4'b00_0_1;
			default :{NS,nSTART,nDOIT} = 4'b00_0_0;
		endcase
	/*****************************************************************/
	//Generate BTU
	/*****************************************************************/
	assign btu_comp = START ? k_half : k;
	assign BTU = btu_comp == Q; 
	
	always @ (*)
		case({DOIT,BTU})
			2'b00: D = 19'b0;
			2'b01: D = 19'b0;
			2'b10: D = Q + 19'b1;
			2'b11: D = 19'b0;
			default: D = 19'b0;
		endcase
	always @(posedge clk, posedge rst)
		if(rst)
			Q <= 19'b0;
		else 
			Q <= D;
			
	/*****************************************************************/
	//Generate DONE
	/*****************************************************************/		
	assign DONE = done_comp == Q1;
	
	always @ (*)
		case({eight,pen})
			2'b00: done_comp = 4'd9;
			2'b01: done_comp = 4'd10;
			2'b10: done_comp = 4'd10;
			2'b11: done_comp = 4'd11;
			default: done_comp = 4'd9;
		endcase
		
	always @ (*)
		case({DOIT,BTU})
			2'b00: D1 = 4'b0;
			2'b01: D1 = 4'b0;
			2'b10: D1 = Q1;
			2'b11: D1 = Q1 + 4'b1;
			default: D1 = 4'b0;
		endcase
	always @ (posedge clk, posedge rst)
		if(rst)
			Q1 <= 4'b0;
		else
			Q1 <= D1;
			
	
	///////////////////////////////////////////////////////////////////
	/////////////////////RECEIVE ENGINE DATA PATH//////////////////////
	///////////////////////////////////////////////////////////////////
	reg [9:0] sr_data, remap_out;
	/*****************************************************************/
	//Shift reg
	/*****************************************************************/		
	assign SH = BTU & (~START);
	
	always @ (posedge clk, posedge rst)
		if(rst)
			sr_data <= 10'b0;
		else 
			if(SH)
				sr_data <= {RX, sr_data[9:1]};
			else 
				sr_data <= sr_data; 
					
	/*****************************************************************/
	//Remap - Combo 
	/*****************************************************************/
	always @(*)
		case ({eight,pen})
			2'b00: remap_out = {2'b00,sr_data[9:2]};
			2'b01: remap_out = {1'b0,sr_data[9:1]};
			2'b10: remap_out = {1'b0,sr_data[9:1]};
			2'b11: remap_out = sr_data;
			default: remap_out = 10'b0;
		endcase 
	/*****************************************************************/
	//RXRDY
	/*****************************************************************/					  
	rs_flop	rxrdy_flop(.clk(clk),
							  .rst(rst),
							  .r(read[0]),
							  .s(DONE),
							  .Q(rxrdy));		

	/*****************************************************************/
	//PERR
	/*****************************************************************/	
	wire par_bit_sel, par_gen_sel, gen_par, perr_set, even, parity; 
	assign even = ohel == 1'b0;
	
	assign par_gen_sel = eight ? remap_out[7] : 1'b0;
	assign par_bit_sel = eight ? remap_out[8] : remap_out[7] ;
	assign parity = par_gen_sel ^ (^remap_out[6:0]);
	assign gen_par = even ? parity : ~parity;
	
	assign perr_set = pen & DONE & (par_bit_sel ^ gen_par); 
	
	rs_flop	perr_flop (.clk(clk),
							  .rst(rst),
							  .r(read[0]),
							  .s(perr_set),
							  .Q(PERR));
	/*****************************************************************/
	//FERR
	/*****************************************************************/	
	wire  ferr_set; 
	reg   st_sel;
	assign ferr_set = DONE & (~st_sel);
	always @ (*)
		case ({eight,pen})
			2'b00: st_sel = remap_out[7];
			2'b01: st_sel = remap_out[8];
			2'b10: st_sel = remap_out[8];
			2'b11: st_sel = remap_out[9];
		endcase	
		
	rs_flop	ferr_flop (.clk(clk),
							  .rst(rst),
							  .r(read[0]),
							  .s(ferr_set),
							  .Q(FERR));
	/*****************************************************************/
	//OVF
	/*****************************************************************/	
	wire ovf_set;
	assign ovf_set = DONE & rxrdy; 
	rs_flop	ovf_flop  (.clk(clk),
							  .rst(rst),
							  .r(read[0]),
							  .s(ovf_set),
							  .Q(OVF));
endmodule
